-- --------------------------------------------------------------------------------
-- Company : Rochester Institute of Technology (RIT )
-- Engineer : Rohan Patil (rnp5285@rit.edu)
--
-- Create Date : 2/19/19
-- Design Name : instr_mem
-- Module Name : instr_mem - behavioral
-- Project Name : ex3
-- Target Devices : Basys3
--
-- Description :  memory module which holds all instructions to fetch  
-- --------------------------------------------------------------------------------

library IEEE ;
use IEEE . STD_LOGIC_1164 .ALL ;
use IEEE . STD_LOGIC_UNSIGNED .ALL;
use IEEE . NUMERIC_STD .ALL;

entity instr_mem is
    port (
            addr : in std_logic_vector(27 downto 0);
            dout : out std_logic_vector(31 downto 0)
    );
end instr_mem;

architecture behav of instr_mem is
    type mem_type is array(0 to 1023) of std_logic_vector(31 downto 0); -- 2^10 size array, checking the first 10 bits of addr
    -- arbitrary memory values
    signal mem : mem_type := (
        
        --PART1
        ---------------------------------------------------------
--         setup, i type add
        0 => "00100000001000010000000000000010",    -- add r1,r1,#2 = 2
        4 => "00100000100000100000000000000001",    -- add r2,r4,#1 = 1
         -- no op
        8 => "00100000000000000000000000000000",   
        12 => "00100000000000000000000000000000",   
        16 => "00100000000000000000000000000000",  
        20 => "00100000000000000000000000000000",   
        
        -- r type
        -- r1 = 1, r1 = 2
        24 => "00000000001000100001100000100000",   -- add r3,r1,r2 = 3
        28 => "00000000001000100001100000100100",   -- and = 0
        32 => "00000000001000100001100000011001",   -- mult = 2 
        36 => "00000000001000100001100000100101",   -- or = 3
        40 => "00000000001000100001100000000000",   -- sll = 4
        44 => "00000000001000100001100000000011",   -- sra = 1
        48 => "00000000001000100001100000000010",   -- srl = 1
        52 => "00000000001000100001100000100011",   -- sub = 1
        56 => "00000000001000100001100000100110",   -- xor = 3
        
        -- j type
        60 => "00001000000000000000000011111010",   -- jump to 1000
        1000=>"00001100000000000000000000010000",   -- jump back to 64
        
        -- i type
        64 => "00100000010000110000000000001111",   -- addi r3,r2,#15 = 16
        68 => "00110000010000110000000000001111",   -- andi = 1
        72 => "00110100010000110000000000001111",   -- ori = 15
        76 => "00111000010000110000000000001111",   -- xori = 1
        80 => "00111100010000110000000000001111",
        84 => "10001100010000110000000000001111",
        
        
-----------------------------------------------------------------------

--        "00100000000000000000000000000000",   

--        -- fibonacci sequence
 --1

--00100000001 00001 0000000000000001 --1
--00100000001 00001 0000000000000000
--00100000001000100000000000000010 --2
--00100000001 00001 0000000000000000
--00100000001 00001 0000000000000011 --3
--00100000001 00001 0000000000000000
--00100000001 00001 0000000000000101 --5
--00100000001 00001 0000000000000000
--00100000001 00001 0000000000001000 --8
--00100000001 00001 0000000000000000
--00100000001 00001 0000000000001101 --13
--00100000001 00001 0000000000000000
--00100000001 00001 0000000000010101 --21
--00100000001 00001 0000000000000000
--00100000001 00001 0000000000100010 --34
--00100000001 00001 0000000000000000
--00100000001 00001 0000000000110111 --55
--00100000001 00001 0000000000000000
        
        

--        0 => "00100000000000010000000000000001", -- ADD R1 <- R0 + 0 = 0 
--        4 => "00100000000000100000000000000001", -- ADD R2 <- R0 + 1 = 1

--        8 => "00100000000000000000000000000000",   
--        12 => "00100000000000000000000000000000",   
--        16 => "00100000000000000000000000000000",   
--        20 => "00100000001000010000000000000001",--   2
--        24 => "00100000000000000000000000000000",   
--        28 => "00100000000000000000000000000000", 
--        32 => "00100000000000000000000000000000",   
--        36 => "00100000001000100000000000000010",--3
--        40 => "00100000000000000000000000000000", 

----        --------------------------------------------
--        44 => "00100000000000000000000000000000", -- r1 <- r1 + r2
--        48 => "00100000000000000000000000000000",   
--        52 => "00100000001000010000000000000011", --  5
--        56 => "00100000000000000000000000000000",   
--        60 => "00100000000000000000000000000000",   
--        64 => "00100000000000000000000000000000",   
--        68 => "00100000001000100000000000001000", -- 8
--        72 => "00100000000000000000000000000000",   
--        76 => "00100000000000000000000000000000",   
--        80 => "00100000000000000000000000000000",     
--        84 => "00100000001000010000000000001101", -- 13
--        88 => "00100000000000000000000000000000", -- jump to 8
--        92 => "00100000000000000000000000000000",
--        96 => "00100000000000000000000000000000",
--        100 => "00100000001000100000000000010101", --21
--        104 => "00100000000000000000000000000000",
--        108 => "00100000000000000000000000000000",
--        112 => "00100000000000000000000000000000",
--        116 => "00100000001000010000000000100010",--
--        120 => "00100000000000000000000000000000",
--        124 => "00100000000000000000000000000000",
--        128 => "00100000000000000000000000000000",
--        132 => "00100000001000100000000000110111", --
--        136 => "00100000000000000000000000000000",
--        140 => "00100000000000000000000000000000",
        
        -- 7 noops
--        0 => "00100000000000010000000000000001", -- ADD R1 <- R0 + 0 = 0 
--        4 => "00100000000000100000000000000001", -- ADD R2 <- R0 + 1 = 1
--        8 => "00100000000000000000000000000000",
--        12 => "00100000000000000000000000000000",
--        16 => "00100000000000000000000000000000",
--        20 => "00100000001000100001000000100000",
--        24 => "00100000000000000000000000000000",
--        28 => "00100000000000000000000000000000",
--        32 => "00100000000000000000000000000000",
--        36 => "00100000000000000000000000000000",
--        40 => "00001000000000000000000000000010", -- JUMP to 8
        
        
        -- no op
--        8 => "00000000000000000000000000000000",   
--        12 => "00000000000000000000000000100000",   
--        16 => "00000000000000000000000000100000",   

        
----        24 => "00000000001000100001100000100000",
--        36 => "00000000000000000000000000100000",
--        40 => "00000000000000000000000000100000",
--        44 => "00000000000000000000000000100000",
--        48 => "00000000000000000000000000100000",
        
--        52 => "00000000001000100010000000100000", -- ADD R3 <- R1+R2
--        56 => "00000000001000100001100000100000",
--        60 => "00000000001000100001100000100000",
--        64 => "00000000001000100001100000100000",
--        68 => "00000000001000100001100000100000",
--        72 => "00000000001000100001100000100000",
--        76 => "00000000001000100001100000100000",
--        80 => "00000000001000100001100000100000",
--        84 => "00000000001000100001100000100000",
--        88 => "00000000001000100001100000100000",
--        92 => "00000000001000100001100000100000",




--        24 => "00000000000000000000000000100000",   
--        28 => "00000000000000000000000000100000",
--        32 => "00000000000000000000000000100000",
        
--        36 => "00000000001000100001100000100000", -- ADD R3 <- R1+R2
--        40 => "00000000000000000000000000100000",   
--        44 => "00000000000000000000000000100000",
--        48 => "00000000000000000000000000100000",
        
--        52 => "00000000010000110010000000100000", -- ADD R4 <- R2+R3
--        56 => "00000000000000000000000000100000",   
--        60 => "00000000000000000000000000100000",
--        64 => "00000000000000000000000000100000",  
            
--        68 => "00000000011001000010100000100000", -- ADD R5 <- R3+R4
--        72 => "00000000000000000000000000100000",   
--        76 => "00000000000000000000000000100000",
--        80 => "00000000000000000000000000100000",
        
--        84 => "00000000100001010011000000100000", -- ADD R6 <- R4+R5
--        88 => "00000000000000000000000000100000",   
--        92 => "00000000000000000000000000100000",
--        96 => "00000000000000000000000000100000",
        
--        100 => "00000000101001100011100000100000", -- ADD R7 <- R5 + R6
--        104 => "00000000000000000000000000100000",   
--        108 => "00000000000000000000000000100000",
--        112 => "00000000000000000000000000100000",
        
        
--        116 => "00000000110001110100000000100000", -- ADD R8 <- R6 + R7
--        120 => "00000000000000000000000000100000",   
--        124 => "00000000000000000000000000100000",
--        128 => "00000000000000000000000000100000",
        
--        132 => "00000000111010000100100000100000", -- ADD R9 <- R7 + R8
--        136 => "00000000000000000000000000100000",   
--        140 => "00000000000000000000000000100000",
--        144 => "00000000000000000000000000100000",
        
--        148 => "00000001000010010101000000100000",  -- ADD R10 <- R8 + R9
--        152 => "00000000000000000000000000100000",   
--        156 => "00000000000000000000000000100000",
--        160 => "00000000000000000000000000100000",


        others=>x"00000000"); -- initialize memory location array
begin
    dout <= mem(to_integer(unsigned(addr(9 downto 0))));    -- dout assigned addr idx of mem
end behav;